library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.numeric_std.ALL;

entity DataMemory is 
	Port (
			Address : in std_logic_vector(31 downto 0);
			WriteData : in std_logic_vector(31 downto 0);
			MemWrite, MemRead : in std_logic;
			ReadData : out std_logic_vector(31 downto 0)
		);
end DataMemory;

architecture Behavioral of DataMemory is

type Memory is array (0 to 30) of std_logic_vector (31 downto 0);  

signal memorySig: Memory:=(
							"00000000000000000000000000000000",	--0
							"00000000000000000000000000000001",	--1 
							"00000000000000000000000000000010",	--2
							"00000000000000000000000000000011",	--3
							"00000000000000000000000000000100",	--4
							"00000000000000000000000000000101",	--5
							"00000000000000000000000000000011",	--6
							"00000000000000000000000000000101",	--7
							"00000000010000110000100000100100",	--8
							"00000000010000110000100000100101",	--9
							"00000000010000110010000000100100",	--10
							"10001100010000010000000000000101",	--11
							"10101100010000010000000000000101",	--12
							"00000000001000000000000101001000",	--13
							"00010100001000100000000000000101",	--14
							"00010100001000100000000000000101",	--15
							"00000000000000000000000000000000",	--16
							"00000000000000000000000000000000",	--17
							"00000000000000000000000000000000",	--18
							"00000000000000000000000000000101",	--19
							"00000000000000000000000000001010",	--20
							"00000000000000000000000000010100",	--21
							"00000000000000000000000000011001",	--22
							"00000000000000000000000000000000",	--23
							"00000000010000110000100000100100",	--24
							"00000000000000000000000000000000",	--25
							"00000000010000110010000000100100",	--26
							"10001100010000010000000000000101",	--27
							"10101100010000010000000000000101",	--28
							"00000000001000000000000101001000",	--29
							"00010100001000100000000000000101"	--30
						);


begin
	
	process(MemWrite,MemRead, Address, WriteData)
	begin
		if(MemWrite='1') then
			memorySig(to_integer(unsigned(Address))) <= WriteData;
		end if;
		if(MemRead='1') then
			ReadData<=memorySig(to_integer(unsigned(Address)));
		end if;
	end process;
	
end Behavioral;
